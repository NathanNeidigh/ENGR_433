module blank ();
endmodule
